`include "awb/provides/heat_transfer_common.bsh"
typedef Bit#(64) CYCLE_COUNTER;

typedef `HEAT_TRANSFER_X_MAX_POINTS N_X_MAX_POINTS;
typedef `HEAT_TRANSFER_Y_MAX_POINTS N_Y_MAX_POINTS;
typedef `HEAT_TRANSFER_X_ENGINE N_X_ENGINES;
typedef `HEAT_TRANSFER_Y_ENGINE N_Y_ENGINES;
typedef TMul#(N_X_ENGINES, N_Y_ENGINES) N_TOTAL_ENGINES;

typedef `HEAT_TRANSFER_NUM_PARTITIONS N_PARTITIONS;
typedef TDiv#(N_TOTAL_ENGINES, N_PARTITIONS) N_ENGINES_PER_PARTITION;

typedef N_ENGINES_PER_PARTITION N_LOCAL_ENGINES;
typedef TMul#(N_ENGINES_PER_PARTITION, n) REMOTE_START_ENGINE#(numeric type n);

typedef TMul#(N_X_MAX_POINTS, N_Y_MAX_POINTS)  N_TOTAL_MAX_POINTS;
typedef Bit#(TAdd#(TAdd#(TLog#(N_X_MAX_POINTS),TLog#(N_Y_MAX_POINTS)),2)) MEM_ADDRESS;
typedef Bit#(`HEAT_TRANSFER_DATA_SIZE) TEST_DATA;

