//----------------------------------------------------------------------//
// The MIT License 
// 
// Copyright (c) 2009 MIT
// 
// Permission is hereby granted, free of charge, to any person 
// obtaining a copy of this software and associated documentation 
// files (the "Software"), to deal in the Software without 
// restriction, including without limitation the rights to use,
// copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
// OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
// HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
// WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
// OTHER DEALINGS IN THE SOFTWARE.
//
// Author: Muralidaran Vijayaraghavan
//
//----------------------------------------------------------------------//

import Types::*;
import List::*;
import Vector::*;
import FixedPointNew::*;

function TData getInverse(Index n);
    Vector#(1000, TData) tempV = Vector::toVector(
            List::cons(0,
            List::cons(fromRational(1,1),
            List::cons(fromRational(1,2),
            List::cons(fromRational(1,3),
            List::cons(fromRational(1,4),
            List::cons(fromRational(1,5),
            List::cons(fromRational(1,6),
            List::cons(fromRational(1,7),
            List::cons(fromRational(1,8),
            List::cons(fromRational(1,9),
            List::cons(fromRational(1,10),
            List::cons(fromRational(1,11),
            List::cons(fromRational(1,12),
            List::cons(fromRational(1,13),
            List::cons(fromRational(1,14),
            List::cons(fromRational(1,15),
            List::cons(fromRational(1,16),
            List::cons(fromRational(1,17),
            List::cons(fromRational(1,18),
            List::cons(fromRational(1,19),
            List::cons(fromRational(1,20),
            List::cons(fromRational(1,21),
            List::cons(fromRational(1,22),
            List::cons(fromRational(1,23),
            List::cons(fromRational(1,24),
            List::cons(fromRational(1,25),
            List::cons(fromRational(1,26),
            List::cons(fromRational(1,27),
            List::cons(fromRational(1,28),
            List::cons(fromRational(1,29),
            List::cons(fromRational(1,30),
            List::cons(fromRational(1,31),
            List::cons(fromRational(1,32),
            List::cons(fromRational(1,33),
            List::cons(fromRational(1,34),
            List::cons(fromRational(1,35),
            List::cons(fromRational(1,36),
            List::cons(fromRational(1,37),
            List::cons(fromRational(1,38),
            List::cons(fromRational(1,39),
            List::cons(fromRational(1,40),
            List::cons(fromRational(1,41),
            List::cons(fromRational(1,42),
            List::cons(fromRational(1,43),
            List::cons(fromRational(1,44),
            List::cons(fromRational(1,45),
            List::cons(fromRational(1,46),
            List::cons(fromRational(1,47),
            List::cons(fromRational(1,48),
            List::cons(fromRational(1,49),
            List::cons(fromRational(1,50),
            List::cons(fromRational(1,51),
            List::cons(fromRational(1,52),
            List::cons(fromRational(1,53),
            List::cons(fromRational(1,54),
            List::cons(fromRational(1,55),
            List::cons(fromRational(1,56),
            List::cons(fromRational(1,57),
            List::cons(fromRational(1,58),
            List::cons(fromRational(1,59),
            List::cons(fromRational(1,60),
            List::cons(fromRational(1,61),
            List::cons(fromRational(1,62),
            List::cons(fromRational(1,63),
            List::cons(fromRational(1,64),
            List::cons(fromRational(1,65),
            List::cons(fromRational(1,66),
            List::cons(fromRational(1,67),
            List::cons(fromRational(1,68),
            List::cons(fromRational(1,69),
            List::cons(fromRational(1,70),
            List::cons(fromRational(1,71),
            List::cons(fromRational(1,72),
            List::cons(fromRational(1,73),
            List::cons(fromRational(1,74),
            List::cons(fromRational(1,75),
            List::cons(fromRational(1,76),
            List::cons(fromRational(1,77),
            List::cons(fromRational(1,78),
            List::cons(fromRational(1,79),
            List::cons(fromRational(1,80),
            List::cons(fromRational(1,81),
            List::cons(fromRational(1,82),
            List::cons(fromRational(1,83),
            List::cons(fromRational(1,84),
            List::cons(fromRational(1,85),
            List::cons(fromRational(1,86),
            List::cons(fromRational(1,87),
            List::cons(fromRational(1,88),
            List::cons(fromRational(1,89),
            List::cons(fromRational(1,90),
            List::cons(fromRational(1,91),
            List::cons(fromRational(1,92),
            List::cons(fromRational(1,93),
            List::cons(fromRational(1,94),
            List::cons(fromRational(1,95),
            List::cons(fromRational(1,96),
            List::cons(fromRational(1,97),
            List::cons(fromRational(1,98),
            List::cons(fromRational(1,99),
            List::cons(fromRational(1,100),
            List::cons(fromRational(1,101),
            List::cons(fromRational(1,102),
            List::cons(fromRational(1,103),
            List::cons(fromRational(1,104),
            List::cons(fromRational(1,105),
            List::cons(fromRational(1,106),
            List::cons(fromRational(1,107),
            List::cons(fromRational(1,108),
            List::cons(fromRational(1,109),
            List::cons(fromRational(1,110),
            List::cons(fromRational(1,111),
            List::cons(fromRational(1,112),
            List::cons(fromRational(1,113),
            List::cons(fromRational(1,114),
            List::cons(fromRational(1,115),
            List::cons(fromRational(1,116),
            List::cons(fromRational(1,117),
            List::cons(fromRational(1,118),
            List::cons(fromRational(1,119),
            List::cons(fromRational(1,120),
            List::cons(fromRational(1,121),
            List::cons(fromRational(1,122),
            List::cons(fromRational(1,123),
            List::cons(fromRational(1,124),
            List::cons(fromRational(1,125),
            List::cons(fromRational(1,126),
            List::cons(fromRational(1,127),
            List::cons(fromRational(1,128),
            List::cons(fromRational(1,129),
            List::cons(fromRational(1,130),
            List::cons(fromRational(1,131),
            List::cons(fromRational(1,132),
            List::cons(fromRational(1,133),
            List::cons(fromRational(1,134),
            List::cons(fromRational(1,135),
            List::cons(fromRational(1,136),
            List::cons(fromRational(1,137),
            List::cons(fromRational(1,138),
            List::cons(fromRational(1,139),
            List::cons(fromRational(1,140),
            List::cons(fromRational(1,141),
            List::cons(fromRational(1,142),
            List::cons(fromRational(1,143),
            List::cons(fromRational(1,144),
            List::cons(fromRational(1,145),
            List::cons(fromRational(1,146),
            List::cons(fromRational(1,147),
            List::cons(fromRational(1,148),
            List::cons(fromRational(1,149),
            List::cons(fromRational(1,150),
            List::cons(fromRational(1,151),
            List::cons(fromRational(1,152),
            List::cons(fromRational(1,153),
            List::cons(fromRational(1,154),
            List::cons(fromRational(1,155),
            List::cons(fromRational(1,156),
            List::cons(fromRational(1,157),
            List::cons(fromRational(1,158),
            List::cons(fromRational(1,159),
            List::cons(fromRational(1,160),
            List::cons(fromRational(1,161),
            List::cons(fromRational(1,162),
            List::cons(fromRational(1,163),
            List::cons(fromRational(1,164),
            List::cons(fromRational(1,165),
            List::cons(fromRational(1,166),
            List::cons(fromRational(1,167),
            List::cons(fromRational(1,168),
            List::cons(fromRational(1,169),
            List::cons(fromRational(1,170),
            List::cons(fromRational(1,171),
            List::cons(fromRational(1,172),
            List::cons(fromRational(1,173),
            List::cons(fromRational(1,174),
            List::cons(fromRational(1,175),
            List::cons(fromRational(1,176),
            List::cons(fromRational(1,177),
            List::cons(fromRational(1,178),
            List::cons(fromRational(1,179),
            List::cons(fromRational(1,180),
            List::cons(fromRational(1,181),
            List::cons(fromRational(1,182),
            List::cons(fromRational(1,183),
            List::cons(fromRational(1,184),
            List::cons(fromRational(1,185),
            List::cons(fromRational(1,186),
            List::cons(fromRational(1,187),
            List::cons(fromRational(1,188),
            List::cons(fromRational(1,189),
            List::cons(fromRational(1,190),
            List::cons(fromRational(1,191),
            List::cons(fromRational(1,192),
            List::cons(fromRational(1,193),
            List::cons(fromRational(1,194),
            List::cons(fromRational(1,195),
            List::cons(fromRational(1,196),
            List::cons(fromRational(1,197),
            List::cons(fromRational(1,198),
            List::cons(fromRational(1,199),
            List::cons(fromRational(1,200),
            List::cons(fromRational(1,201),
            List::cons(fromRational(1,202),
            List::cons(fromRational(1,203),
            List::cons(fromRational(1,204),
            List::cons(fromRational(1,205),
            List::cons(fromRational(1,206),
            List::cons(fromRational(1,207),
            List::cons(fromRational(1,208),
            List::cons(fromRational(1,209),
            List::cons(fromRational(1,210),
            List::cons(fromRational(1,211),
            List::cons(fromRational(1,212),
            List::cons(fromRational(1,213),
            List::cons(fromRational(1,214),
            List::cons(fromRational(1,215),
            List::cons(fromRational(1,216),
            List::cons(fromRational(1,217),
            List::cons(fromRational(1,218),
            List::cons(fromRational(1,219),
            List::cons(fromRational(1,220),
            List::cons(fromRational(1,221),
            List::cons(fromRational(1,222),
            List::cons(fromRational(1,223),
            List::cons(fromRational(1,224),
            List::cons(fromRational(1,225),
            List::cons(fromRational(1,226),
            List::cons(fromRational(1,227),
            List::cons(fromRational(1,228),
            List::cons(fromRational(1,229),
            List::cons(fromRational(1,230),
            List::cons(fromRational(1,231),
            List::cons(fromRational(1,232),
            List::cons(fromRational(1,233),
            List::cons(fromRational(1,234),
            List::cons(fromRational(1,235),
            List::cons(fromRational(1,236),
            List::cons(fromRational(1,237),
            List::cons(fromRational(1,238),
            List::cons(fromRational(1,239),
            List::cons(fromRational(1,240),
            List::cons(fromRational(1,241),
            List::cons(fromRational(1,242),
            List::cons(fromRational(1,243),
            List::cons(fromRational(1,244),
            List::cons(fromRational(1,245),
            List::cons(fromRational(1,246),
            List::cons(fromRational(1,247),
            List::cons(fromRational(1,248),
            List::cons(fromRational(1,249),
            List::cons(fromRational(1,250),
            List::cons(fromRational(1,251),
            List::cons(fromRational(1,252),
            List::cons(fromRational(1,253),
            List::cons(fromRational(1,254),
            List::cons(fromRational(1,255),
            List::cons(fromRational(1,256),
            List::cons(fromRational(1,257),
            List::cons(fromRational(1,258),
            List::cons(fromRational(1,259),
            List::cons(fromRational(1,260),
            List::cons(fromRational(1,261),
            List::cons(fromRational(1,262),
            List::cons(fromRational(1,263),
            List::cons(fromRational(1,264),
            List::cons(fromRational(1,265),
            List::cons(fromRational(1,266),
            List::cons(fromRational(1,267),
            List::cons(fromRational(1,268),
            List::cons(fromRational(1,269),
            List::cons(fromRational(1,270),
            List::cons(fromRational(1,271),
            List::cons(fromRational(1,272),
            List::cons(fromRational(1,273),
            List::cons(fromRational(1,274),
            List::cons(fromRational(1,275),
            List::cons(fromRational(1,276),
            List::cons(fromRational(1,277),
            List::cons(fromRational(1,278),
            List::cons(fromRational(1,279),
            List::cons(fromRational(1,280),
            List::cons(fromRational(1,281),
            List::cons(fromRational(1,282),
            List::cons(fromRational(1,283),
            List::cons(fromRational(1,284),
            List::cons(fromRational(1,285),
            List::cons(fromRational(1,286),
            List::cons(fromRational(1,287),
            List::cons(fromRational(1,288),
            List::cons(fromRational(1,289),
            List::cons(fromRational(1,290),
            List::cons(fromRational(1,291),
            List::cons(fromRational(1,292),
            List::cons(fromRational(1,293),
            List::cons(fromRational(1,294),
            List::cons(fromRational(1,295),
            List::cons(fromRational(1,296),
            List::cons(fromRational(1,297),
            List::cons(fromRational(1,298),
            List::cons(fromRational(1,299),
            List::cons(fromRational(1,300),
            List::cons(fromRational(1,301),
            List::cons(fromRational(1,302),
            List::cons(fromRational(1,303),
            List::cons(fromRational(1,304),
            List::cons(fromRational(1,305),
            List::cons(fromRational(1,306),
            List::cons(fromRational(1,307),
            List::cons(fromRational(1,308),
            List::cons(fromRational(1,309),
            List::cons(fromRational(1,310),
            List::cons(fromRational(1,311),
            List::cons(fromRational(1,312),
            List::cons(fromRational(1,313),
            List::cons(fromRational(1,314),
            List::cons(fromRational(1,315),
            List::cons(fromRational(1,316),
            List::cons(fromRational(1,317),
            List::cons(fromRational(1,318),
            List::cons(fromRational(1,319),
            List::cons(fromRational(1,320),
            List::cons(fromRational(1,321),
            List::cons(fromRational(1,322),
            List::cons(fromRational(1,323),
            List::cons(fromRational(1,324),
            List::cons(fromRational(1,325),
            List::cons(fromRational(1,326),
            List::cons(fromRational(1,327),
            List::cons(fromRational(1,328),
            List::cons(fromRational(1,329),
            List::cons(fromRational(1,330),
            List::cons(fromRational(1,331),
            List::cons(fromRational(1,332),
            List::cons(fromRational(1,333),
            List::cons(fromRational(1,334),
            List::cons(fromRational(1,335),
            List::cons(fromRational(1,336),
            List::cons(fromRational(1,337),
            List::cons(fromRational(1,338),
            List::cons(fromRational(1,339),
            List::cons(fromRational(1,340),
            List::cons(fromRational(1,341),
            List::cons(fromRational(1,342),
            List::cons(fromRational(1,343),
            List::cons(fromRational(1,344),
            List::cons(fromRational(1,345),
            List::cons(fromRational(1,346),
            List::cons(fromRational(1,347),
            List::cons(fromRational(1,348),
            List::cons(fromRational(1,349),
            List::cons(fromRational(1,350),
            List::cons(fromRational(1,351),
            List::cons(fromRational(1,352),
            List::cons(fromRational(1,353),
            List::cons(fromRational(1,354),
            List::cons(fromRational(1,355),
            List::cons(fromRational(1,356),
            List::cons(fromRational(1,357),
            List::cons(fromRational(1,358),
            List::cons(fromRational(1,359),
            List::cons(fromRational(1,360),
            List::cons(fromRational(1,361),
            List::cons(fromRational(1,362),
            List::cons(fromRational(1,363),
            List::cons(fromRational(1,364),
            List::cons(fromRational(1,365),
            List::cons(fromRational(1,366),
            List::cons(fromRational(1,367),
            List::cons(fromRational(1,368),
            List::cons(fromRational(1,369),
            List::cons(fromRational(1,370),
            List::cons(fromRational(1,371),
            List::cons(fromRational(1,372),
            List::cons(fromRational(1,373),
            List::cons(fromRational(1,374),
            List::cons(fromRational(1,375),
            List::cons(fromRational(1,376),
            List::cons(fromRational(1,377),
            List::cons(fromRational(1,378),
            List::cons(fromRational(1,379),
            List::cons(fromRational(1,380),
            List::cons(fromRational(1,381),
            List::cons(fromRational(1,382),
            List::cons(fromRational(1,383),
            List::cons(fromRational(1,384),
            List::cons(fromRational(1,385),
            List::cons(fromRational(1,386),
            List::cons(fromRational(1,387),
            List::cons(fromRational(1,388),
            List::cons(fromRational(1,389),
            List::cons(fromRational(1,390),
            List::cons(fromRational(1,391),
            List::cons(fromRational(1,392),
            List::cons(fromRational(1,393),
            List::cons(fromRational(1,394),
            List::cons(fromRational(1,395),
            List::cons(fromRational(1,396),
            List::cons(fromRational(1,397),
            List::cons(fromRational(1,398),
            List::cons(fromRational(1,399),
            List::cons(fromRational(1,400),
            List::cons(fromRational(1,401),
            List::cons(fromRational(1,402),
            List::cons(fromRational(1,403),
            List::cons(fromRational(1,404),
            List::cons(fromRational(1,405),
            List::cons(fromRational(1,406),
            List::cons(fromRational(1,407),
            List::cons(fromRational(1,408),
            List::cons(fromRational(1,409),
            List::cons(fromRational(1,410),
            List::cons(fromRational(1,411),
            List::cons(fromRational(1,412),
            List::cons(fromRational(1,413),
            List::cons(fromRational(1,414),
            List::cons(fromRational(1,415),
            List::cons(fromRational(1,416),
            List::cons(fromRational(1,417),
            List::cons(fromRational(1,418),
            List::cons(fromRational(1,419),
            List::cons(fromRational(1,420),
            List::cons(fromRational(1,421),
            List::cons(fromRational(1,422),
            List::cons(fromRational(1,423),
            List::cons(fromRational(1,424),
            List::cons(fromRational(1,425),
            List::cons(fromRational(1,426),
            List::cons(fromRational(1,427),
            List::cons(fromRational(1,428),
            List::cons(fromRational(1,429),
            List::cons(fromRational(1,430),
            List::cons(fromRational(1,431),
            List::cons(fromRational(1,432),
            List::cons(fromRational(1,433),
            List::cons(fromRational(1,434),
            List::cons(fromRational(1,435),
            List::cons(fromRational(1,436),
            List::cons(fromRational(1,437),
            List::cons(fromRational(1,438),
            List::cons(fromRational(1,439),
            List::cons(fromRational(1,440),
            List::cons(fromRational(1,441),
            List::cons(fromRational(1,442),
            List::cons(fromRational(1,443),
            List::cons(fromRational(1,444),
            List::cons(fromRational(1,445),
            List::cons(fromRational(1,446),
            List::cons(fromRational(1,447),
            List::cons(fromRational(1,448),
            List::cons(fromRational(1,449),
            List::cons(fromRational(1,450),
            List::cons(fromRational(1,451),
            List::cons(fromRational(1,452),
            List::cons(fromRational(1,453),
            List::cons(fromRational(1,454),
            List::cons(fromRational(1,455),
            List::cons(fromRational(1,456),
            List::cons(fromRational(1,457),
            List::cons(fromRational(1,458),
            List::cons(fromRational(1,459),
            List::cons(fromRational(1,460),
            List::cons(fromRational(1,461),
            List::cons(fromRational(1,462),
            List::cons(fromRational(1,463),
            List::cons(fromRational(1,464),
            List::cons(fromRational(1,465),
            List::cons(fromRational(1,466),
            List::cons(fromRational(1,467),
            List::cons(fromRational(1,468),
            List::cons(fromRational(1,469),
            List::cons(fromRational(1,470),
            List::cons(fromRational(1,471),
            List::cons(fromRational(1,472),
            List::cons(fromRational(1,473),
            List::cons(fromRational(1,474),
            List::cons(fromRational(1,475),
            List::cons(fromRational(1,476),
            List::cons(fromRational(1,477),
            List::cons(fromRational(1,478),
            List::cons(fromRational(1,479),
            List::cons(fromRational(1,480),
            List::cons(fromRational(1,481),
            List::cons(fromRational(1,482),
            List::cons(fromRational(1,483),
            List::cons(fromRational(1,484),
            List::cons(fromRational(1,485),
            List::cons(fromRational(1,486),
            List::cons(fromRational(1,487),
            List::cons(fromRational(1,488),
            List::cons(fromRational(1,489),
            List::cons(fromRational(1,490),
            List::cons(fromRational(1,491),
            List::cons(fromRational(1,492),
            List::cons(fromRational(1,493),
            List::cons(fromRational(1,494),
            List::cons(fromRational(1,495),
            List::cons(fromRational(1,496),
            List::cons(fromRational(1,497),
            List::cons(fromRational(1,498),
            List::cons(fromRational(1,499),
            List::cons(fromRational(1,500),
            List::cons(fromRational(1,501),
            List::cons(fromRational(1,502),
            List::cons(fromRational(1,503),
            List::cons(fromRational(1,504),
            List::cons(fromRational(1,505),
            List::cons(fromRational(1,506),
            List::cons(fromRational(1,507),
            List::cons(fromRational(1,508),
            List::cons(fromRational(1,509),
            List::cons(fromRational(1,510),
            List::cons(fromRational(1,511),
            List::cons(fromRational(1,512),
            List::cons(fromRational(1,513),
            List::cons(fromRational(1,514),
            List::cons(fromRational(1,515),
            List::cons(fromRational(1,516),
            List::cons(fromRational(1,517),
            List::cons(fromRational(1,518),
            List::cons(fromRational(1,519),
            List::cons(fromRational(1,520),
            List::cons(fromRational(1,521),
            List::cons(fromRational(1,522),
            List::cons(fromRational(1,523),
            List::cons(fromRational(1,524),
            List::cons(fromRational(1,525),
            List::cons(fromRational(1,526),
            List::cons(fromRational(1,527),
            List::cons(fromRational(1,528),
            List::cons(fromRational(1,529),
            List::cons(fromRational(1,530),
            List::cons(fromRational(1,531),
            List::cons(fromRational(1,532),
            List::cons(fromRational(1,533),
            List::cons(fromRational(1,534),
            List::cons(fromRational(1,535),
            List::cons(fromRational(1,536),
            List::cons(fromRational(1,537),
            List::cons(fromRational(1,538),
            List::cons(fromRational(1,539),
            List::cons(fromRational(1,540),
            List::cons(fromRational(1,541),
            List::cons(fromRational(1,542),
            List::cons(fromRational(1,543),
            List::cons(fromRational(1,544),
            List::cons(fromRational(1,545),
            List::cons(fromRational(1,546),
            List::cons(fromRational(1,547),
            List::cons(fromRational(1,548),
            List::cons(fromRational(1,549),
            List::cons(fromRational(1,550),
            List::cons(fromRational(1,551),
            List::cons(fromRational(1,552),
            List::cons(fromRational(1,553),
            List::cons(fromRational(1,554),
            List::cons(fromRational(1,555),
            List::cons(fromRational(1,556),
            List::cons(fromRational(1,557),
            List::cons(fromRational(1,558),
            List::cons(fromRational(1,559),
            List::cons(fromRational(1,560),
            List::cons(fromRational(1,561),
            List::cons(fromRational(1,562),
            List::cons(fromRational(1,563),
            List::cons(fromRational(1,564),
            List::cons(fromRational(1,565),
            List::cons(fromRational(1,566),
            List::cons(fromRational(1,567),
            List::cons(fromRational(1,568),
            List::cons(fromRational(1,569),
            List::cons(fromRational(1,570),
            List::cons(fromRational(1,571),
            List::cons(fromRational(1,572),
            List::cons(fromRational(1,573),
            List::cons(fromRational(1,574),
            List::cons(fromRational(1,575),
            List::cons(fromRational(1,576),
            List::cons(fromRational(1,577),
            List::cons(fromRational(1,578),
            List::cons(fromRational(1,579),
            List::cons(fromRational(1,580),
            List::cons(fromRational(1,581),
            List::cons(fromRational(1,582),
            List::cons(fromRational(1,583),
            List::cons(fromRational(1,584),
            List::cons(fromRational(1,585),
            List::cons(fromRational(1,586),
            List::cons(fromRational(1,587),
            List::cons(fromRational(1,588),
            List::cons(fromRational(1,589),
            List::cons(fromRational(1,590),
            List::cons(fromRational(1,591),
            List::cons(fromRational(1,592),
            List::cons(fromRational(1,593),
            List::cons(fromRational(1,594),
            List::cons(fromRational(1,595),
            List::cons(fromRational(1,596),
            List::cons(fromRational(1,597),
            List::cons(fromRational(1,598),
            List::cons(fromRational(1,599),
            List::cons(fromRational(1,600),
            List::cons(fromRational(1,601),
            List::cons(fromRational(1,602),
            List::cons(fromRational(1,603),
            List::cons(fromRational(1,604),
            List::cons(fromRational(1,605),
            List::cons(fromRational(1,606),
            List::cons(fromRational(1,607),
            List::cons(fromRational(1,608),
            List::cons(fromRational(1,609),
            List::cons(fromRational(1,610),
            List::cons(fromRational(1,611),
            List::cons(fromRational(1,612),
            List::cons(fromRational(1,613),
            List::cons(fromRational(1,614),
            List::cons(fromRational(1,615),
            List::cons(fromRational(1,616),
            List::cons(fromRational(1,617),
            List::cons(fromRational(1,618),
            List::cons(fromRational(1,619),
            List::cons(fromRational(1,620),
            List::cons(fromRational(1,621),
            List::cons(fromRational(1,622),
            List::cons(fromRational(1,623),
            List::cons(fromRational(1,624),
            List::cons(fromRational(1,625),
            List::cons(fromRational(1,626),
            List::cons(fromRational(1,627),
            List::cons(fromRational(1,628),
            List::cons(fromRational(1,629),
            List::cons(fromRational(1,630),
            List::cons(fromRational(1,631),
            List::cons(fromRational(1,632),
            List::cons(fromRational(1,633),
            List::cons(fromRational(1,634),
            List::cons(fromRational(1,635),
            List::cons(fromRational(1,636),
            List::cons(fromRational(1,637),
            List::cons(fromRational(1,638),
            List::cons(fromRational(1,639),
            List::cons(fromRational(1,640),
            List::cons(fromRational(1,641),
            List::cons(fromRational(1,642),
            List::cons(fromRational(1,643),
            List::cons(fromRational(1,644),
            List::cons(fromRational(1,645),
            List::cons(fromRational(1,646),
            List::cons(fromRational(1,647),
            List::cons(fromRational(1,648),
            List::cons(fromRational(1,649),
            List::cons(fromRational(1,650),
            List::cons(fromRational(1,651),
            List::cons(fromRational(1,652),
            List::cons(fromRational(1,653),
            List::cons(fromRational(1,654),
            List::cons(fromRational(1,655),
            List::cons(fromRational(1,656),
            List::cons(fromRational(1,657),
            List::cons(fromRational(1,658),
            List::cons(fromRational(1,659),
            List::cons(fromRational(1,660),
            List::cons(fromRational(1,661),
            List::cons(fromRational(1,662),
            List::cons(fromRational(1,663),
            List::cons(fromRational(1,664),
            List::cons(fromRational(1,665),
            List::cons(fromRational(1,666),
            List::cons(fromRational(1,667),
            List::cons(fromRational(1,668),
            List::cons(fromRational(1,669),
            List::cons(fromRational(1,670),
            List::cons(fromRational(1,671),
            List::cons(fromRational(1,672),
            List::cons(fromRational(1,673),
            List::cons(fromRational(1,674),
            List::cons(fromRational(1,675),
            List::cons(fromRational(1,676),
            List::cons(fromRational(1,677),
            List::cons(fromRational(1,678),
            List::cons(fromRational(1,679),
            List::cons(fromRational(1,680),
            List::cons(fromRational(1,681),
            List::cons(fromRational(1,682),
            List::cons(fromRational(1,683),
            List::cons(fromRational(1,684),
            List::cons(fromRational(1,685),
            List::cons(fromRational(1,686),
            List::cons(fromRational(1,687),
            List::cons(fromRational(1,688),
            List::cons(fromRational(1,689),
            List::cons(fromRational(1,690),
            List::cons(fromRational(1,691),
            List::cons(fromRational(1,692),
            List::cons(fromRational(1,693),
            List::cons(fromRational(1,694),
            List::cons(fromRational(1,695),
            List::cons(fromRational(1,696),
            List::cons(fromRational(1,697),
            List::cons(fromRational(1,698),
            List::cons(fromRational(1,699),
            List::cons(fromRational(1,700),
            List::cons(fromRational(1,701),
            List::cons(fromRational(1,702),
            List::cons(fromRational(1,703),
            List::cons(fromRational(1,704),
            List::cons(fromRational(1,705),
            List::cons(fromRational(1,706),
            List::cons(fromRational(1,707),
            List::cons(fromRational(1,708),
            List::cons(fromRational(1,709),
            List::cons(fromRational(1,710),
            List::cons(fromRational(1,711),
            List::cons(fromRational(1,712),
            List::cons(fromRational(1,713),
            List::cons(fromRational(1,714),
            List::cons(fromRational(1,715),
            List::cons(fromRational(1,716),
            List::cons(fromRational(1,717),
            List::cons(fromRational(1,718),
            List::cons(fromRational(1,719),
            List::cons(fromRational(1,720),
            List::cons(fromRational(1,721),
            List::cons(fromRational(1,722),
            List::cons(fromRational(1,723),
            List::cons(fromRational(1,724),
            List::cons(fromRational(1,725),
            List::cons(fromRational(1,726),
            List::cons(fromRational(1,727),
            List::cons(fromRational(1,728),
            List::cons(fromRational(1,729),
            List::cons(fromRational(1,730),
            List::cons(fromRational(1,731),
            List::cons(fromRational(1,732),
            List::cons(fromRational(1,733),
            List::cons(fromRational(1,734),
            List::cons(fromRational(1,735),
            List::cons(fromRational(1,736),
            List::cons(fromRational(1,737),
            List::cons(fromRational(1,738),
            List::cons(fromRational(1,739),
            List::cons(fromRational(1,740),
            List::cons(fromRational(1,741),
            List::cons(fromRational(1,742),
            List::cons(fromRational(1,743),
            List::cons(fromRational(1,744),
            List::cons(fromRational(1,745),
            List::cons(fromRational(1,746),
            List::cons(fromRational(1,747),
            List::cons(fromRational(1,748),
            List::cons(fromRational(1,749),
            List::cons(fromRational(1,750),
            List::cons(fromRational(1,751),
            List::cons(fromRational(1,752),
            List::cons(fromRational(1,753),
            List::cons(fromRational(1,754),
            List::cons(fromRational(1,755),
            List::cons(fromRational(1,756),
            List::cons(fromRational(1,757),
            List::cons(fromRational(1,758),
            List::cons(fromRational(1,759),
            List::cons(fromRational(1,760),
            List::cons(fromRational(1,761),
            List::cons(fromRational(1,762),
            List::cons(fromRational(1,763),
            List::cons(fromRational(1,764),
            List::cons(fromRational(1,765),
            List::cons(fromRational(1,766),
            List::cons(fromRational(1,767),
            List::cons(fromRational(1,768),
            List::cons(fromRational(1,769),
            List::cons(fromRational(1,770),
            List::cons(fromRational(1,771),
            List::cons(fromRational(1,772),
            List::cons(fromRational(1,773),
            List::cons(fromRational(1,774),
            List::cons(fromRational(1,775),
            List::cons(fromRational(1,776),
            List::cons(fromRational(1,777),
            List::cons(fromRational(1,778),
            List::cons(fromRational(1,779),
            List::cons(fromRational(1,780),
            List::cons(fromRational(1,781),
            List::cons(fromRational(1,782),
            List::cons(fromRational(1,783),
            List::cons(fromRational(1,784),
            List::cons(fromRational(1,785),
            List::cons(fromRational(1,786),
            List::cons(fromRational(1,787),
            List::cons(fromRational(1,788),
            List::cons(fromRational(1,789),
            List::cons(fromRational(1,790),
            List::cons(fromRational(1,791),
            List::cons(fromRational(1,792),
            List::cons(fromRational(1,793),
            List::cons(fromRational(1,794),
            List::cons(fromRational(1,795),
            List::cons(fromRational(1,796),
            List::cons(fromRational(1,797),
            List::cons(fromRational(1,798),
            List::cons(fromRational(1,799),
            List::cons(fromRational(1,800),
            List::cons(fromRational(1,801),
            List::cons(fromRational(1,802),
            List::cons(fromRational(1,803),
            List::cons(fromRational(1,804),
            List::cons(fromRational(1,805),
            List::cons(fromRational(1,806),
            List::cons(fromRational(1,807),
            List::cons(fromRational(1,808),
            List::cons(fromRational(1,809),
            List::cons(fromRational(1,810),
            List::cons(fromRational(1,811),
            List::cons(fromRational(1,812),
            List::cons(fromRational(1,813),
            List::cons(fromRational(1,814),
            List::cons(fromRational(1,815),
            List::cons(fromRational(1,816),
            List::cons(fromRational(1,817),
            List::cons(fromRational(1,818),
            List::cons(fromRational(1,819),
            List::cons(fromRational(1,820),
            List::cons(fromRational(1,821),
            List::cons(fromRational(1,822),
            List::cons(fromRational(1,823),
            List::cons(fromRational(1,824),
            List::cons(fromRational(1,825),
            List::cons(fromRational(1,826),
            List::cons(fromRational(1,827),
            List::cons(fromRational(1,828),
            List::cons(fromRational(1,829),
            List::cons(fromRational(1,830),
            List::cons(fromRational(1,831),
            List::cons(fromRational(1,832),
            List::cons(fromRational(1,833),
            List::cons(fromRational(1,834),
            List::cons(fromRational(1,835),
            List::cons(fromRational(1,836),
            List::cons(fromRational(1,837),
            List::cons(fromRational(1,838),
            List::cons(fromRational(1,839),
            List::cons(fromRational(1,840),
            List::cons(fromRational(1,841),
            List::cons(fromRational(1,842),
            List::cons(fromRational(1,843),
            List::cons(fromRational(1,844),
            List::cons(fromRational(1,845),
            List::cons(fromRational(1,846),
            List::cons(fromRational(1,847),
            List::cons(fromRational(1,848),
            List::cons(fromRational(1,849),
            List::cons(fromRational(1,850),
            List::cons(fromRational(1,851),
            List::cons(fromRational(1,852),
            List::cons(fromRational(1,853),
            List::cons(fromRational(1,854),
            List::cons(fromRational(1,855),
            List::cons(fromRational(1,856),
            List::cons(fromRational(1,857),
            List::cons(fromRational(1,858),
            List::cons(fromRational(1,859),
            List::cons(fromRational(1,860),
            List::cons(fromRational(1,861),
            List::cons(fromRational(1,862),
            List::cons(fromRational(1,863),
            List::cons(fromRational(1,864),
            List::cons(fromRational(1,865),
            List::cons(fromRational(1,866),
            List::cons(fromRational(1,867),
            List::cons(fromRational(1,868),
            List::cons(fromRational(1,869),
            List::cons(fromRational(1,870),
            List::cons(fromRational(1,871),
            List::cons(fromRational(1,872),
            List::cons(fromRational(1,873),
            List::cons(fromRational(1,874),
            List::cons(fromRational(1,875),
            List::cons(fromRational(1,876),
            List::cons(fromRational(1,877),
            List::cons(fromRational(1,878),
            List::cons(fromRational(1,879),
            List::cons(fromRational(1,880),
            List::cons(fromRational(1,881),
            List::cons(fromRational(1,882),
            List::cons(fromRational(1,883),
            List::cons(fromRational(1,884),
            List::cons(fromRational(1,885),
            List::cons(fromRational(1,886),
            List::cons(fromRational(1,887),
            List::cons(fromRational(1,888),
            List::cons(fromRational(1,889),
            List::cons(fromRational(1,890),
            List::cons(fromRational(1,891),
            List::cons(fromRational(1,892),
            List::cons(fromRational(1,893),
            List::cons(fromRational(1,894),
            List::cons(fromRational(1,895),
            List::cons(fromRational(1,896),
            List::cons(fromRational(1,897),
            List::cons(fromRational(1,898),
            List::cons(fromRational(1,899),
            List::cons(fromRational(1,900),
            List::cons(fromRational(1,901),
            List::cons(fromRational(1,902),
            List::cons(fromRational(1,903),
            List::cons(fromRational(1,904),
            List::cons(fromRational(1,905),
            List::cons(fromRational(1,906),
            List::cons(fromRational(1,907),
            List::cons(fromRational(1,908),
            List::cons(fromRational(1,909),
            List::cons(fromRational(1,910),
            List::cons(fromRational(1,911),
            List::cons(fromRational(1,912),
            List::cons(fromRational(1,913),
            List::cons(fromRational(1,914),
            List::cons(fromRational(1,915),
            List::cons(fromRational(1,916),
            List::cons(fromRational(1,917),
            List::cons(fromRational(1,918),
            List::cons(fromRational(1,919),
            List::cons(fromRational(1,920),
            List::cons(fromRational(1,921),
            List::cons(fromRational(1,922),
            List::cons(fromRational(1,923),
            List::cons(fromRational(1,924),
            List::cons(fromRational(1,925),
            List::cons(fromRational(1,926),
            List::cons(fromRational(1,927),
            List::cons(fromRational(1,928),
            List::cons(fromRational(1,929),
            List::cons(fromRational(1,930),
            List::cons(fromRational(1,931),
            List::cons(fromRational(1,932),
            List::cons(fromRational(1,933),
            List::cons(fromRational(1,934),
            List::cons(fromRational(1,935),
            List::cons(fromRational(1,936),
            List::cons(fromRational(1,937),
            List::cons(fromRational(1,938),
            List::cons(fromRational(1,939),
            List::cons(fromRational(1,940),
            List::cons(fromRational(1,941),
            List::cons(fromRational(1,942),
            List::cons(fromRational(1,943),
            List::cons(fromRational(1,944),
            List::cons(fromRational(1,945),
            List::cons(fromRational(1,946),
            List::cons(fromRational(1,947),
            List::cons(fromRational(1,948),
            List::cons(fromRational(1,949),
            List::cons(fromRational(1,950),
            List::cons(fromRational(1,951),
            List::cons(fromRational(1,952),
            List::cons(fromRational(1,953),
            List::cons(fromRational(1,954),
            List::cons(fromRational(1,955),
            List::cons(fromRational(1,956),
            List::cons(fromRational(1,957),
            List::cons(fromRational(1,958),
            List::cons(fromRational(1,959),
            List::cons(fromRational(1,960),
            List::cons(fromRational(1,961),
            List::cons(fromRational(1,962),
            List::cons(fromRational(1,963),
            List::cons(fromRational(1,964),
            List::cons(fromRational(1,965),
            List::cons(fromRational(1,966),
            List::cons(fromRational(1,967),
            List::cons(fromRational(1,968),
            List::cons(fromRational(1,969),
            List::cons(fromRational(1,970),
            List::cons(fromRational(1,971),
            List::cons(fromRational(1,972),
            List::cons(fromRational(1,973),
            List::cons(fromRational(1,974),
            List::cons(fromRational(1,975),
            List::cons(fromRational(1,976),
            List::cons(fromRational(1,977),
            List::cons(fromRational(1,978),
            List::cons(fromRational(1,979),
            List::cons(fromRational(1,980),
            List::cons(fromRational(1,981),
            List::cons(fromRational(1,982),
            List::cons(fromRational(1,983),
            List::cons(fromRational(1,984),
            List::cons(fromRational(1,985),
            List::cons(fromRational(1,986),
            List::cons(fromRational(1,987),
            List::cons(fromRational(1,988),
            List::cons(fromRational(1,989),
            List::cons(fromRational(1,990),
            List::cons(fromRational(1,991),
            List::cons(fromRational(1,992),
            List::cons(fromRational(1,993),
            List::cons(fromRational(1,994),
            List::cons(fromRational(1,995),
            List::cons(fromRational(1,996),
            List::cons(fromRational(1,997),
            List::cons(fromRational(1,998),
            List::cons(fromRational(1,999),
   List::nil)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
   return tempV[n];
endfunction
